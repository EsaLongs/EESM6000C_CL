`define ADDER_SIZE 128
`define MUL_SIZE 64

// You can set MUL_SIZE as 8, 16, 32, 64, 128 ....
// But you must make sure ADDER_SIZE = 2 * MUL_SIZE