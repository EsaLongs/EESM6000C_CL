module booth4multiplier_onestage (
  ports
);
  
endmodule