//---------------------- Original Code -----------------------//
