//---------------------- Original Code -----------------------//
  //---------------------- Code 1 ----------------------------//
  if (condition) begin
    foo = bar;
  end 
  else begin
    foo = bum;
  end

  //---------------------- Code 2 ----------------------------//
  assign a=((addr&mask)==My_addr)?b[1]:!b[0];

  //---------------------- Code 3 ----------------------------//
  logic [7:0][3:0] data[128] [2];

  //---------------------- Code 4 ----------------------------//
  typedef logic[31:0]word_t;

  //---------------------- Code 5 ----------------------------//
  assign foo = condition_a ? condition_a_x ? x : y : b;

//---------------------- Modified Code -----------------------//
  //---------------------- Code 1 ----------------------------//
  // End else begin must be together on one line
  if (condition) begin
    foo = bar;
  end else begin
    foo = bum;
  end

  //---------------------- Code 2 ----------------------------//
  // Include whitespace on both sides of all binary operators
  assign a = ((addr & mask) == My_addr) ? b[1] : !b[0];

  //---------------------- Code 3 ----------------------------//
  // There must not be a space between dimensions
  logic [7:0][3:0] data[128][2];

  //---------------------- Code 4 ----------------------------//
  // There must be a space around packed dimensions
  typedef logic [31:0] word_t;

  //---------------------- Code 5 ----------------------------//
  // Ternary expressions nested in the true condition of another ternary expression must be enclosed in parentheses
  assign foo = condition_a ? (condition_a_x ? x : y) : b;