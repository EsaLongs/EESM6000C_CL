module moduleName (
  ports
);
  
endmodule