module moduleName #(
  parameter  = ;

) (
  ports
);
  
endmodule