module brent_kung_adder (
  ports
);
endmodule