`define ADDER_SIZE 64