/*
In order to satisfy all the flip-flops timing requirement, 
which both paths should have a delay under 10, we need to 
adjust some of the combinational logic part in path#2 and 
put them in path#1. The ideal situation is both of them 
have a delay of 9.

*/