//---------------------- Original Code -----------------------//