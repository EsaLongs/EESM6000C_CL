`define ADDER_SIZE 32