`define ADDER_SIZE 64 // Can be ste as 16 * n